/*
 * Copyright (c) 2025. All rights reserved.
 * Created by enrique, 17/05/25
 */

class Transaction;

    function automatic new ();

    endfunction : new

    virtual function automatic void display (string name);

    endfunction : display
endclass : Transaction